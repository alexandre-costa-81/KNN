library ieee;
package example_type is
    type example_float32 is array(0 to 74) of STD_LOGIC_VECTOR(31 DOWNTO 0);
end package example_type;

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_SIGNED.all;
use IEEE.math_real.all;
use ieee.numeric_std.all;
use work.example_type.all;
--------------------------------------

entity test_receive is

port(
	CLOCK_50: in std_logic;
	UART_TXD: OUT STD_LOGIC;
	UART_RXD: IN STD_LOGIC;
	KEY: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	LEDR: OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
	LEDG: OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
);
end test_receive;

architecture KNN_arch of test_receive is
type example75f is array(0 to 74) of std_logic_vector(31 downto 0);
type examples is array(0 to 1) of example75f;
signal x: example75f;
signal exemplos: examples;
signal starting: std_logic := '1';
signal temp_r: float32;
signal minDist: float32:="01111111011111111111111111111111";
SIGNAL TX_DATA: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL TX_START: STD_LOGIC := '0';
SIGNAL TX_BUSY: STD_LOGIC;
SIGNAL RX_DATA: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL RX_BUSY: STD_LOGIC;
SIGNAL WORD_INDEX: INTEGER RANGE 0 TO 3:=0;
SIGNAL DATA0: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL DATA1: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL DATA2: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL DATA3: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL COLUMN: INTEGER RANGE 0 TO 74:=0;
SIGNAL receiving: integer range 0 to 3 := 0;
COMPONENT TX
PORT(
CLK: IN STD_LOGIC;
START: IN STD_LOGIC;
BUSY: OUT STD_LOGIC;
DATA: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
TX_LINE: OUT STD_LOGIC
);
END COMPONENT TX;
COMPONENT RX
PORT(
CLK: IN STD_LOGIC;
RX_LINE: IN STD_LOGIC;
DATA: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
BUSY: OUT STD_LOGIC
);
END COMPONENT RX;
BEGIN
	C1: TX PORT MAP(CLOCK_50, TX_START, TX_BUSY, TX_DATA, UART_TXD);
	C2: RX PORT MAP(CLOCK_50, UART_RXD, RX_DATA, RX_BUSY);  
	PROCESS(CLOCK_50)
	variable y: std_logic;
	variable etapa: integer range 0 to 10:=0;
	variable countc: integer range 0 to 77:=0;
	variable countr: integer range 0 to 77:=0;
	variable count_wait: integer range 0 to 5000002:=0;
	BEGIN	
		IF(CLOCK_50'EVENT AND CLOCK_50='1') THEN
			IF(receiving=0 AND TX_BUSY='0') THEN
				TX_DATA <= "11111111";
				TX_START <= '1';
				receiving <= 1;
			ELSE
				TX_START <= '0';
			END IF;
			IF(receiving = 1 AND RX_BUSY='0') THEN
				IF(WORD_INDEX=0) THEN
					DATA0 <= RX_DATA;
					WORD_INDEX <= WORD_INDEX+1;
				ELSIF(WORD_INDEX=1) THEN
					DATA1 <= RX_DATA;
					WORD_INDEX <= WORD_INDEX+1;
				ELSIF(WORD_INDEX=2) THEN
					DATA2 <= RX_DATA;
					WORD_INDEX <= WORD_INDEX+1;
				ELSIF(WORD_INDEX=3) THEN
					DATA3 <= RX_DATA;
					x(COLUMN) <= DATA0 & DATA1 & DATA2 & DATA3;
					COLUMN <= COLUMN + 1;
					WORD_INDEX <= 0;
					IF(COLUMN = 75) THEN --75, 0 to 74
						COLUMN <= 0;
						--LEDR(17 DOWNTO 0) <= x(2)(17 DOWNTO 0);
						receiving <= 2;
					END IF;
				END IF;
			end if;
			--Calculate KNN and display result
			if(receiving = 2) then
				if(etapa = 0) then
					--if key is pressed, each time, of 2 times, could record example frame, class 1, then class 2
					--better to use one switch, when '0', on next loop, get first example, then when '1', get next example
					--if(SW(0)='0') then
					--	receiving <= 2;
					--end if;
					if(starting = '1') then
						--example of arm up(one class), and down(other class)
						exemplos <= ((
"00111101100100110011101010001010",
"00111111000100100100011100000010",
"00111111110110011110001111000001",
"00111101101001011101111100100010",
"00111110110101101101001010001001",
"00111111110110010110010111000011",
"00111101101000111011010011110110",
"00111110101100001100011000101110",
"00111111110110000011100011000001",
"00111101100111000000000110100011",
"00111101111010100101100111000000",
"00111111110100111000001101101011",
"00111110011110111111010100001110",
"00111110100001010100110011011011",
"00111111110100101001000101100100",
"10111101110110110011111100100001",
"00111110100010111110110111111010",
"00111111110101001100101001001111",
"00111101100011111101010000111001",
"10111110010100110111010100000000",
"00111111110010111100000011011011",
"00111110000101110111100000010100",
"10111110010011101010000101000000",
"00111111110001101001000010011011",
"10111100001100010010110100110100",
"10111110010011100101010100111011",
"00111111110001110101100001100100",
"00111110101000101010111010001110",
"00111100010010011000111001010100",
"00111111110011011000011100000101",
"00111110101100110001101100010101",
"10111110001111101111110001111010",
"00111111110000101010100101110001",
"00111110101011001010000011000011",
"10111110011001000001100111100011",
"00111111110000000011101000111011",
"00111110101010110110101000011111",
"10111110100100010001101010111001",
"00111111101111001111111111100011",
"00111110100111000011001001100110",
"10111110011001000001101101110110",
"00111111101111100010000011100110",
"10111110001011000000010101001111",
"00111101000011010000001101010011",
"00111111110011001010000010001000",
"10111110010010100110110000011010",
"10111110001000001100100101010100",
"00111111101111110101010001100101",
"10111110001111111010001101110111",
"10111110001010010100011100000110",
"00111111101111111000100010110001",
"10111110001110101011100010100110",
"10111110011010000011011000100010",
"00111111101111001100010111001010",
"10111101111100100001011110001111",
"10111110001111111101000111011101",
"00111111110000111111011101001001",
"00111110001011100001000100010010",
"10111111000010101000100101010101",
"00111111110000010100000111011001",
"00111110001001110000111110111111",
"10111111011100110101100100110110",
"00111111110001001101011100111000",
"00111110000111110010010100011100",
"10111111011101101001101101001010",
"00111111101100100001111010011011",
"10111101010100100101001101010100",
"10111111000010011111001111111001",
"00111111110000000010001111001000",
"10111101100110001100000010001011",
"10111111011100101111110110010111",
"00111111110000100111011000001000",
"10111101100111101010110101001111",
"10111111011101100011000111010111",
"00111111101011111011110100111000"),
(
"10111011110111010001111001010100",
"00111111000100110111101100111001",
"00111111110110101000000010110110",
"10111011100000101000001111010011",
"00111110110110111010100010000010",
"00111111110110001101111001100101",
"10111000001101000101101011100110",
"00111110101101100101000010000011",
"00111111110101111110101000001100",
"00111100010001110000110010011001",
"00111110000001000111110011111010",
"00111111110100111101111111000010",
"00111110010001110110010100110100",
"00111110100110011000101001000100",
"00111111110100110011101101011100",
"10111110010011010001100100010101",
"00111110100101011010111100101001",
"00111111110100101111101111111100",
"00111100111011100110110110011100",
"10111110001111100110000010000000",
"00111111110011010000100100011000",
"00111101110111101000000000111001",
"10111110001101111100011000110010",
"00111111110010001001010111101010",
"10111101010101000011000001101110",
"10111110001111000000101101010110",
"00111111110001111101110101011101",
"00111110110000110010001100110110",
"00111110101001110111100010011010",
"00111111110001000011100000010001",
"00111110110011011011111001111111",
"00111111000010110101111010010110",
"00111111101111001011001001111101",
"00111110110100110100111010111010",
"00111111001001010010101001100011",
"00111111101111001000111010100100",
"00111110110100111010011110111001",
"00111111001101111010111111001001",
"00111111101110100110111100100110",
"00111110111010100111000010001111",
"00111111000111110101101101100000",
"00111111101110111000111110110100",
"10111110110000111111101110011100",
"00111110101110010111101011101110",
"00111111110001000100001001011011",
"10111110110100101111101001110010",
"00111111000100010110011110001000",
"00111111101110011101000111001100",
"10111110110100010011011000011110",
"00111111001010001011001011011001",
"00111111101110100110011101000001",
"10111110110101001001010011010101",
"00111111001111001011001100011100",
"00111111101110010011001010000011",
"10111110111010001001000011110111",
"00111111001010001000100010100100",
"00111111101110000101010110110000",
"00111110001100011011010011111110",
"10111111000000111101000001101100",
"00111111101111110011110110000110",
"00111110010101101111111101111110",
"10111111011010111001100110000000",
"00111111110000011000110011101011",
"00111110010100100011011011000001",
"10111111011011110000111110111111",
"00111111101011101100111111100001",
"10111101101011110110001001110100",
"10111111000001000001111110100111",
"00111111101111101001010011110111",
"10111101011100100001101000101110",
"10111111011011100000000000101010",
"00111111110000010100010110101110",
"10111101011011100111011100001100",
"10111111011100010110001111001100",
"00111111101011101000010101001101"));

						starting <= '0';
					end if;
					minDist <= "01111111011111111111111111111111";
					temp_r <= "00000000000000000000000000000000";
					countc := 0;
					countr := 0;
					etapa := 1;
				elsif(etapa = 1) then --acquire frame from Kinect
					--send byte to start receiving frame, if key is pressed
						--wait for key otherwise
						--or loop. Receive, process, give class. 
						--		Better. 
						--Just leave out key. 
					--IF(KEY(0)='0' AND TX_BUSY='0') THEN --no need, just loop, always ask for example
--					IF(TX_BUSY='0') THEN
--						TX_DATA <= "11111111";
--						TX_START <= '1';
--						receiving <= 1;
--					ELSE
--						TX_START<='0';
--					END IF;
					etapa := 2;
				elsif(etapa = 2) then
					--testo <= to_slv(minDist);
					if(countr = 2) then --rows of example
						count_wait := 0;
						etapa := 3;
					else
						--co <= countc;
						if(countc = 75) then --columns of example
							--check to see if distance is lower
							--temp_b <= temp_r;
							if(temp_r < minDist) then
								minDist <= temp_r;
								if(countr = 0) then
									y := '0';
								else
									y := '1';
								end if;
							end if; 
							countc := countc + 1;
							countr := countr + 1;
							--testo <= to_slv(temp_r);
						elsif(countc = 76) then --columns of example
							--testo <= to_slv(minDist);
							--etapa := 3;
							countc := 0;
							count_wait := 0;
							temp_r <= "00000000000000000000000000000000";
						else
							--cw <= count_wait;
							if(count_wait = 0) then
								--temp_r := temp_r + ((to_float(exemplos(0)(countr)) - to_float(x(countr))) * (to_float(to_float(exemplos(0)(countr)) - to_float(testi_b))));
								--temp_r := temp_r + sqrt((to_float(exemplos(0)(countr)) - to_float(x(countr))) * (to_float(exemplos(0)(countr)) - to_float(x(countr))));				
								temp_r <= temp_r + ((to_float(exemplos(countr)(countc)) - to_float(x(countc))) * (to_float(exemplos(countr)(countc)) - to_float(x(countc))));				
								--temp_r <= to_float(exemplos(countr)(countc));
								--co <= countr;
								count_wait := count_wait + 1;
							elsif(count_wait = 10) then
								countc := countc + 1;
								count_wait := 0;
								--testo <= to_slv(temp_r);
							else
								count_wait := count_wait + 1;
							end if;
						end if;
					end if;
				elsif(etapa = 3) then
					--testo <= to_slv(temp_r);
					--turn on all green or red leds, depending on class
					--yy <= y;
					if(count_wait = 5000000) then
						if(y = '0') then
							LEDR(17 DOWNTO 0) <= (others => '1');
							LEDG(8 DOWNTO 0) <= (others => '0');
						else
							LEDR(17 DOWNTO 0) <= (others => '0');
							LEDG(8 DOWNTO 0) <= (others => '1');
						end if;
						receiving <= 0;
						etapa := 0;
						count_wait := 0;
					else
						count_wait := count_wait + 1;
					end if;
					--go back to start
				end if;
			end if;
		END IF;
	END PROCESS;
end KNN_arch;